module ysyx_220066_cpu(

)

endmodule