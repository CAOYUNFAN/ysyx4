module ysyx_220066_Ex(

)

endmodule

module ysyx_220066_ALU(

)

endmodule

module ysyx_220066_nxtPC(

)

endmodule